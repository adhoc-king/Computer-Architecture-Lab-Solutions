module decoder5_32(register,reg_no);
	input [4:0] reg_no;
	output [31:0] register;
	assign register[0] = (~reg_no[4] & ~reg_no[3] & ~reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[1] = (~reg_no[4] & ~reg_no[3] & ~reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[2] = (~reg_no[4] & ~reg_no[3] & ~reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[3] = (~reg_no[4] & ~reg_no[3] & ~reg_no[2] & reg_no[1] & reg_no[0]),
	    register[4] = (~reg_no[4] & ~reg_no[3] & reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[5] = (~reg_no[4] & ~reg_no[3] & reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[6] = (~reg_no[4] & ~reg_no[3] & reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[7] = (~reg_no[4] & ~reg_no[3] & reg_no[2] & reg_no[1] & reg_no[0]),
	    register[8] = (~reg_no[4] & reg_no[3] & ~reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[9] = (~reg_no[4] & reg_no[3] & ~reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[10] = (~reg_no[4] & reg_no[3] & ~reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[11] = (~reg_no[4] & reg_no[3] & ~reg_no[2] & reg_no[1] & reg_no[0]),
	    register[12] = (~reg_no[4] & reg_no[3] & reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[13] = (~reg_no[4] & reg_no[3] & reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[14] = (~reg_no[4] & reg_no[3] & reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[15] = (~reg_no[4] & reg_no[3] & reg_no[2] & reg_no[1] & reg_no[0]),
	    register[16] = (reg_no[4] & ~reg_no[3] & ~reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[17] = (reg_no[4] & ~reg_no[3] & ~reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[18] = (reg_no[4] & ~reg_no[3] & ~reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[19] = (reg_no[4] & ~reg_no[3] & ~reg_no[2] & reg_no[1] & reg_no[0]),
	    register[20] = (reg_no[4] & ~reg_no[3] & reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[21] = (reg_no[4] & ~reg_no[3] & reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[22] = (reg_no[4] & ~reg_no[3] & reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[23] = (reg_no[4] & ~reg_no[3] & reg_no[2] & reg_no[1] & reg_no[0]),
	    register[24] = (reg_no[4] & reg_no[3] & ~reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[25] = (reg_no[4] & reg_no[3] & ~reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[26] = (reg_no[4] & reg_no[3] & ~reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[27] = (reg_no[4] & reg_no[3] & ~reg_no[2] & reg_no[1] & reg_no[0]),
	    register[28] = (reg_no[4] & reg_no[3] & reg_no[2] & ~reg_no[1] & ~reg_no[0]),
	    register[29] = (reg_no[4] & reg_no[3] & reg_no[2] & ~reg_no[1] & reg_no[0]),
	    register[30] = (reg_no[4] & reg_no[3] & reg_no[2] & reg_no[1] & ~reg_no[0]),
	    register[31] = (reg_no[4] & reg_no[3] & reg_no[2] & reg_no[1] & reg_no[0]);
endmodule 