module Encrypt(cipherText, plainText, key);
	
endmodule