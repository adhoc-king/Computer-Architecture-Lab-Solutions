module mux16to1_test;
	wire out;
	reg [15:0] in;
	reg [3:0] sel;
	mux16to1_gate mux(out, in, sel);
	initial
	begin
		$monitor($time, " out=%b in=%b, sel=%b", out, in, sel);
		#0 in=16'b1000000000000000;
		#3 in=16'b0100000000000000;
		#3 in=16'b0010000000000000;
		#3 in=16'b0001000000000000;
		#3 in=16'b0000100000000000;
		#3 in=16'b0000010000000000;
		#3 in=16'b0000001000000000;
		#3 in=16'b0000000100000000;
		#3 in=16'b0000000010000000;
		#3 in=16'b0000000001000000;
		#3 in=16'b0000000000100000;
		#3 in=16'b0000000000010000;
		#3 in=16'b0000000000001000;
		#3 in=16'b0000000000000100;
		#3 in=16'b0000000000000010;
		#3 in=16'b0000000000000001;
	end
	initial
	begin
		#0 sel = 4'b0000;
		repeat(15) #3 sel = sel + 4'b0001;
	end
endmodule