module InstructionMemory(Instruction, PC, clock);
	input [5:0] PC;
	input clock;
	output [31:0] Instruction;
	reg [31:0] Instruction;
	reg [31:0] Memory [0:31];
	initial
	begin
		Memory[0] = 32'b00000000000000000000000000000000;
		Memory[1] = 32'b00000000000000000000000001010100;
		Memory[2] = 32'b00000000000000000000000000001011;
		Memory[4] = 32'b00000000000000000000000000000000;
		Memory[5] = 32'b00000000000000000000000000000000;
		Memory[6] = 32'b00000000000000000000000000000000;
		Memory[7] = 32'b00000000000000000000000000000000;
		Memory[8] = 32'b00000000000000000000000000000000;
		Memory[9] = 32'b00000000000000000000000000000000;
		Memory[10] = 32'b00000000000000000000000000000000;
		Memory[11] = 32'b00000000000000000000000000000000;
		Memory[12] = 32'b00000000000000000000000000000000;
		Memory[13] = 32'b00000000000000000000000000000000;
		Memory[14] = 32'b00000000000000000000000000000000;
		Memory[15] = 32'b00000000000000000000000000000000;
		Memory[16] = 32'b00000000000000000000000000000000;
		Memory[17] = 32'b00000000000000000000000000000000;
		Memory[18] = 32'b00000000000000000000000000000000;
		Memory[19] = 32'b00000000000000000000000000000000;
		Memory[20] = 32'b00000000000000000000000000000000;
		Memory[21] = 32'b00000000000000000000000000000000;
		Memory[22] = 32'b00000000000000000000000000000000;
		Memory[23] = 32'b00000000000000000000000000000000;
		Memory[24] = 32'b00000000000000000000000000000000;
		Memory[25] = 32'b00000000000000000000000000000000;
		Memory[26] = 32'b00000000000000000000000000000000;
		Memory[27] = 32'b00000000000000000000000000000000;
		Memory[28] = 32'b00000000000000000000000000000000;
		Memory[29] = 32'b00000000000000000000000000000000;
		Memory[30] = 32'b00000000000000000000000000000000;
		Memory[31] = 32'b00000000000000000000000000000000;
	end
	always @(posedge clock)
		Instruction = Memory[PC/4];
endmodule